**.subckt untitled
XM1 __UNCONNECTED_PIN__0 __UNCONNECTED_PIN__1 net1 GND sky130_fd_pr__nfet_05v0_nvt L=0.300 W=0.6 nf=1
+ ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net1 __UNCONNECTED_PIN__2 __UNCONNECTED_PIN__3 GND sky130_fd_pr__nfet_05v0_nvt L=0.15 W=0.175 nf=1
+ ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM3 __UNCONNECTED_PIN__4 __UNCONNECTED_PIN__5 net1 GND sky130_fd_pr__nfet_05v0_nvt L=0.300 W=0.6 nf=1
+ ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
**.ends
** flattened .save nodes
.end
